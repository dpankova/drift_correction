////////////////////////////////////////////////////////////////
// Daria Pankova Wed Jul 22 12:20:07 EDT 2015
// test_rom.v
//
// "Pseudo RAM with baseline data"
// A custom Verilog HDL module.
// 
////////////////////////////////////////////////////////////////


module test_rom_example(
		input [8:0]   rdaddr,
		output [13:0] adc_val 
		);
   reg [13:0] adc_rom[0:511];
   
   assign adc_val = adc_rom[rdaddr];
   
   initial begin
      adc_rom[0] <= 4780;
      adc_rom[1] <= 4779;
      adc_rom[2] <= 4775;
      adc_rom[3] <= 4777;
      adc_rom[4] <= 4775;
      adc_rom[5] <= 4782;
      adc_rom[6] <= 4775;
      adc_rom[7] <= 4777;
      adc_rom[8] <= 4780;
      adc_rom[9] <= 4779;
      adc_rom[10] <= 4779;
      adc_rom[11] <= 4775;
      adc_rom[12] <= 4778;
      adc_rom[13] <= 4780;
      adc_rom[14] <= 4773;
      adc_rom[15] <= 4780;
      adc_rom[16] <= 4780;
      adc_rom[17] <= 4780;
      adc_rom[18] <= 4780;
      adc_rom[19] <= 4775;
      adc_rom[20] <= 4777;
      adc_rom[21] <= 4781;
      adc_rom[22] <= 4776;
      adc_rom[23] <= 4779;
      adc_rom[24] <= 4772;
      adc_rom[25] <= 4781;
      adc_rom[26] <= 4777;
      adc_rom[27] <= 4780;
      adc_rom[28] <= 4778;
      adc_rom[29] <= 4777;
      adc_rom[30] <= 4779;
      adc_rom[31] <= 4779;
      adc_rom[32] <= 4777;
      adc_rom[33] <= 4779;
      adc_rom[34] <= 4773;
      adc_rom[35] <= 4780;
      adc_rom[36] <= 4774;
      adc_rom[37] <= 4775;
      adc_rom[38] <= 4777;
      adc_rom[39] <= 4776;
      adc_rom[40] <= 4774;
      adc_rom[41] <= 4777;
      adc_rom[42] <= 4778;
      adc_rom[43] <= 4778;
      adc_rom[44] <= 4778;
      adc_rom[45] <= 4780;
      adc_rom[46] <= 4774;
      adc_rom[47] <= 4777;
      adc_rom[48] <= 4776;
      adc_rom[49] <= 4778;
      adc_rom[50] <= 4782;
      adc_rom[51] <= 4776;
      adc_rom[52] <= 4776;
      adc_rom[53] <= 4777;
      adc_rom[54] <= 4778;
      adc_rom[55] <= 4778;
      adc_rom[56] <= 4772;
      adc_rom[57] <= 4778;
      adc_rom[58] <= 4777;
      adc_rom[59] <= 4777;
      adc_rom[60] <= 4779;
      adc_rom[61] <= 4776;
      adc_rom[62] <= 4783;
      adc_rom[63] <= 4781;
      adc_rom[64] <= 4772;
      adc_rom[65] <= 4781;
      adc_rom[66] <= 4775;
      adc_rom[67] <= 4776;
      adc_rom[68] <= 4778;
      adc_rom[69] <= 4776;
      adc_rom[70] <= 4773;
      adc_rom[71] <= 4779;
      adc_rom[72] <= 4780;
      adc_rom[73] <= 4779;
      adc_rom[74] <= 4779;
      adc_rom[75] <= 4779;
      adc_rom[76] <= 4778;
      adc_rom[77] <= 4774;
      adc_rom[78] <= 4779;
      adc_rom[79] <= 4770;
      adc_rom[80] <= 4781;
      adc_rom[81] <= 4776;
      adc_rom[82] <= 4779;
      adc_rom[83] <= 4778;
      adc_rom[84] <= 4775;
      adc_rom[85] <= 4777;
      adc_rom[86] <= 4768;
      adc_rom[87] <= 4776;
      adc_rom[88] <= 4776;
      adc_rom[89] <= 4773;
      adc_rom[90] <= 4781;
      adc_rom[91] <= 4774;
      adc_rom[92] <= 4779;
      adc_rom[93] <= 4781;
      adc_rom[94] <= 4772;
      adc_rom[95] <= 4780;
      adc_rom[96] <= 4773;
      adc_rom[97] <= 4775;
      adc_rom[98] <= 4777;
      adc_rom[99] <= 4777;
      adc_rom[100] <= 4783;
      adc_rom[101] <= 4777;
      adc_rom[102] <= 4774;
      adc_rom[103] <= 4780;
      adc_rom[104] <= 4771;
      adc_rom[105] <= 4781;
      adc_rom[106] <= 4778;
      adc_rom[107] <= 4773;
      adc_rom[108] <= 4780;
      adc_rom[109] <= 4780;
      adc_rom[110] <= 4782;
      adc_rom[111] <= 4776;
      adc_rom[112] <= 4778;
      adc_rom[113] <= 4782;
      adc_rom[114] <= 4776;
      adc_rom[115] <= 4785;
      adc_rom[116] <= 4777;
      adc_rom[117] <= 4777;
      adc_rom[118] <= 4776;
      adc_rom[119] <= 4775;
      adc_rom[120] <= 4778;
      adc_rom[121] <= 4774;
      adc_rom[122] <= 4777;
      adc_rom[123] <= 4779;
      adc_rom[124] <= 4777;
      adc_rom[125] <= 4781;
      adc_rom[126] <= 4777;
      adc_rom[127] <= 4778;
      adc_rom[128] <= 4777;
      adc_rom[129] <= 4777;
      adc_rom[130] <= 4779;
      adc_rom[131] <= 4775;
      adc_rom[132] <= 4778;
      adc_rom[133] <= 4779;
      adc_rom[134] <= 4776;
      adc_rom[135] <= 4779;
      adc_rom[136] <= 4778;
      adc_rom[137] <= 4778;
      adc_rom[138] <= 4779;
      adc_rom[139] <= 4775;
      adc_rom[140] <= 4777;
      adc_rom[141] <= 4778;
      adc_rom[142] <= 4777;
      adc_rom[143] <= 4780;
      adc_rom[144] <= 4773;
      adc_rom[145] <= 4781;
      adc_rom[146] <= 4776;
      adc_rom[147] <= 4775;
      adc_rom[148] <= 4775;
      adc_rom[149] <= 4777;
      adc_rom[150] <= 4782;
      adc_rom[151] <= 4776;
      adc_rom[152] <= 4776;
      adc_rom[153] <= 4776;
      adc_rom[154] <= 4774;
      adc_rom[155] <= 4777;
      adc_rom[156] <= 4770;
      adc_rom[157] <= 4776;
      adc_rom[158] <= 4778;
      adc_rom[159] <= 4778;
      adc_rom[160] <= 4778;
      adc_rom[161] <= 4778;
      adc_rom[162] <= 4772;
      adc_rom[163] <= 4778;
      adc_rom[164] <= 4772;
      adc_rom[165] <= 4784;
      adc_rom[166] <= 4775;
      adc_rom[167] <= 4775;
      adc_rom[168] <= 4779;
      adc_rom[169] <= 4779;
      adc_rom[170] <= 4780;
      adc_rom[171] <= 4777;
      adc_rom[172] <= 4777;
      adc_rom[173] <= 4777;
      adc_rom[174] <= 4776;
      adc_rom[175] <= 4781;
      adc_rom[176] <= 4779;
      adc_rom[177] <= 4774;
      adc_rom[178] <= 4779;
      adc_rom[179] <= 4778;
      adc_rom[180] <= 4780;
      adc_rom[181] <= 4776;
      adc_rom[182] <= 4776;
      adc_rom[183] <= 4779;
      adc_rom[184] <= 4776;
      adc_rom[185] <= 4783;
      adc_rom[186] <= 4776;
      adc_rom[187] <= 4774;
      adc_rom[188] <= 4779;
      adc_rom[189] <= 4778;
      adc_rom[190] <= 4782;
      adc_rom[191] <= 4774;
      adc_rom[192] <= 4774;
      adc_rom[193] <= 4781;
      adc_rom[194] <= 4774;
      adc_rom[195] <= 4780;
      adc_rom[196] <= 4773;
      adc_rom[197] <= 4777;
      adc_rom[198] <= 4779;
      adc_rom[199] <= 4774;
      adc_rom[200] <= 4777;
      adc_rom[201] <= 4776;
      adc_rom[202] <= 4777;
      adc_rom[203] <= 4775;
      adc_rom[204] <= 4777;
      adc_rom[205] <= 4777;
      adc_rom[206] <= 4775;
      adc_rom[207] <= 4773;
      adc_rom[208] <= 4779;
      adc_rom[209] <= 4777;
      adc_rom[210] <= 4782;
      adc_rom[211] <= 4775;
      adc_rom[212] <= 4780;
      adc_rom[213] <= 4779;
      adc_rom[214] <= 4773;
      adc_rom[215] <= 4775;
      adc_rom[216] <= 4774;
      adc_rom[217] <= 4772;
      adc_rom[218] <= 4781;
      adc_rom[219] <= 4776;
      adc_rom[220] <= 4773;
      adc_rom[221] <= 4778;
      adc_rom[222] <= 4777;
      adc_rom[223] <= 4781;
      adc_rom[224] <= 4772;
      adc_rom[225] <= 4784;
      adc_rom[226] <= 4777;
      adc_rom[227] <= 4776;
      adc_rom[228] <= 4778;
      adc_rom[229] <= 4775;
      adc_rom[230] <= 4776;
      adc_rom[231] <= 4775;
      adc_rom[232] <= 4779;
      adc_rom[233] <= 4780;
      adc_rom[234] <= 4775;
      adc_rom[235] <= 4783;
      adc_rom[236] <= 4775;
      adc_rom[237] <= 4778;
      adc_rom[238] <= 4779;
      adc_rom[239] <= 4771;
      adc_rom[240] <= 4778;
      adc_rom[241] <= 4779;
      adc_rom[242] <= 4778;
      adc_rom[243] <= 4778;
      adc_rom[244] <= 4775;
      adc_rom[245] <= 4781;
      adc_rom[246] <= 4775;
      adc_rom[247] <= 4779;
      adc_rom[248] <= 4777;
      adc_rom[249] <= 4774;
      adc_rom[250] <= 4781;
      adc_rom[251] <= 4777;
      adc_rom[252] <= 4779;
      adc_rom[253] <= 4781;
      adc_rom[254] <= 4777;
      adc_rom[255] <= 4779;
      adc_rom[256] <= 4778;
      adc_rom[257] <= 4777;
      adc_rom[258] <= 4774;
      adc_rom[259] <= 4774;
      adc_rom[260] <= 4780;
      adc_rom[261] <= 4780;
      adc_rom[262] <= 4778;
      adc_rom[263] <= 4778;
      adc_rom[264] <= 4772;
      adc_rom[265] <= 4781;
      adc_rom[266] <= 4776;
      adc_rom[267] <= 4779;
      adc_rom[268] <= 4775;
      adc_rom[269] <= 4776;
      adc_rom[270] <= 4783;
      adc_rom[271] <= 4771;
      adc_rom[272] <= 4776;
      adc_rom[273] <= 4784;
      adc_rom[274] <= 4773;
      adc_rom[275] <= 4783;
      adc_rom[276] <= 4771;
      adc_rom[277] <= 4782;
      adc_rom[278] <= 4779;
      adc_rom[279] <= 4774;
      adc_rom[280] <= 4776;
      adc_rom[281] <= 4773;
      adc_rom[282] <= 4779;
      adc_rom[283] <= 4780;
      adc_rom[284] <= 4773;
      adc_rom[285] <= 4777;
      adc_rom[286] <= 4780;
      adc_rom[287] <= 4776;
      adc_rom[288] <= 4773;
      adc_rom[289] <= 4780;
      adc_rom[290] <= 4779;
      adc_rom[291] <= 4774;
      adc_rom[292] <= 4772;
      adc_rom[293] <= 4777;
      adc_rom[294] <= 4775;
      adc_rom[295] <= 4774;
      adc_rom[296] <= 4772;
      adc_rom[297] <= 4776;
      adc_rom[298] <= 4780;
      adc_rom[299] <= 4776;
      adc_rom[300] <= 4774;
      adc_rom[301] <= 4776;
      adc_rom[302] <= 4779;
      adc_rom[303] <= 4774;
      adc_rom[304] <= 4773;
      adc_rom[305] <= 4780;
      adc_rom[306] <= 4775;
      adc_rom[307] <= 4774;
      adc_rom[308] <= 4778;
      adc_rom[309] <= 4772;
      adc_rom[310] <= 4779;
      adc_rom[311] <= 4777;
      adc_rom[312] <= 4774;
      adc_rom[313] <= 4777;
      adc_rom[314] <= 4775;
      adc_rom[315] <= 4781;
      adc_rom[316] <= 4774;
      adc_rom[317] <= 4779;
      adc_rom[318] <= 4779;
      adc_rom[319] <= 4774;
      adc_rom[320] <= 4777;
      adc_rom[321] <= 4778;
      adc_rom[322] <= 4779;
      adc_rom[323] <= 4775;
      adc_rom[324] <= 4776;
      adc_rom[325] <= 4780;
      adc_rom[326] <= 4778;
      adc_rom[327] <= 4774;
      adc_rom[328] <= 4783;
      adc_rom[329] <= 4775;
      adc_rom[330] <= 4781;
      adc_rom[331] <= 4776;
      adc_rom[332] <= 4777;
      adc_rom[333] <= 4782;
      adc_rom[334] <= 4776;
      adc_rom[335] <= 4781;
      adc_rom[336] <= 4776;
      adc_rom[337] <= 4775;
      adc_rom[338] <= 4783;
      adc_rom[339] <= 4773;
      adc_rom[340] <= 4776;
      adc_rom[341] <= 4772;
      adc_rom[342] <= 4773;
      adc_rom[343] <= 4778;
      adc_rom[344] <= 4771;
      adc_rom[345] <= 4780;
      adc_rom[346] <= 4776;
      adc_rom[347] <= 4772;
      adc_rom[348] <= 4778;
      adc_rom[349] <= 4776;
      adc_rom[350] <= 4780;
      adc_rom[351] <= 4773;
      adc_rom[352] <= 4776;
      adc_rom[353] <= 4776;
      adc_rom[354] <= 4775;
      adc_rom[355] <= 4777;
      adc_rom[356] <= 4775;
      adc_rom[357] <= 4775;
      adc_rom[358] <= 4780;
      adc_rom[359] <= 4775;
      adc_rom[360] <= 4780;
      adc_rom[361] <= 4775;
      adc_rom[362] <= 4776;
      adc_rom[363] <= 4778;
      adc_rom[364] <= 4775;
      adc_rom[365] <= 4778;
      adc_rom[366] <= 4776;
      adc_rom[367] <= 4775;
      adc_rom[368] <= 4774;
      adc_rom[369] <= 4776;
      adc_rom[370] <= 4782;
      adc_rom[371] <= 4770;
      adc_rom[372] <= 4775;
      adc_rom[373] <= 4777;
      adc_rom[374] <= 4774;
      adc_rom[375] <= 4778;
      adc_rom[376] <= 4775;
      adc_rom[377] <= 4776;
      adc_rom[378] <= 4777;
      adc_rom[379] <= 4772;
      adc_rom[380] <= 4775;
      adc_rom[381] <= 4775;
      adc_rom[382] <= 4777;
      adc_rom[383] <= 4779;
      adc_rom[384] <= 4774;
      adc_rom[385] <= 4780;
      adc_rom[386] <= 4779;
      adc_rom[387] <= 4777;
      adc_rom[388] <= 4779;
      adc_rom[389] <= 4778;
      adc_rom[390] <= 4777;
      adc_rom[391] <= 4776;
      adc_rom[392] <= 4775;
      adc_rom[393] <= 4782;
      adc_rom[394] <= 4773;
      adc_rom[395] <= 4780;
      adc_rom[396] <= 4774;
      adc_rom[397] <= 4781;
      adc_rom[398] <= 4774;
      adc_rom[399] <= 4782;
      adc_rom[400] <= 4775;
      adc_rom[401] <= 4774;
      adc_rom[402] <= 4780;
      adc_rom[403] <= 4779;
      adc_rom[404] <= 4777;
      adc_rom[405] <= 4782;
      adc_rom[406] <= 4772;
      adc_rom[407] <= 4778;
      adc_rom[408] <= 4772;
      adc_rom[409] <= 4773;
      adc_rom[410] <= 4785;
      adc_rom[411] <= 4772;
      adc_rom[412] <= 4779;
      adc_rom[413] <= 4780;
      adc_rom[414] <= 4768;
      adc_rom[415] <= 4777;
      adc_rom[416] <= 4778;
      adc_rom[417] <= 4779;
      adc_rom[418] <= 4780;
      adc_rom[419] <= 4776;
      adc_rom[420] <= 4778;
      adc_rom[421] <= 4779;
      adc_rom[422] <= 4773;
      adc_rom[423] <= 4784;
      adc_rom[424] <= 4773;
      adc_rom[425] <= 4779;
      adc_rom[426] <= 4777;
      adc_rom[427] <= 4779;
      adc_rom[428] <= 4775;
      adc_rom[429] <= 4774;
      adc_rom[430] <= 4780;
      adc_rom[431] <= 4776;
      adc_rom[432] <= 4773;
      adc_rom[433] <= 4776;
      adc_rom[434] <= 4771;
      adc_rom[435] <= 4777;
      adc_rom[436] <= 4774;
      adc_rom[437] <= 4775;
      adc_rom[438] <= 4778;
      adc_rom[439] <= 4775;
      adc_rom[440] <= 4780;
      adc_rom[441] <= 4775;
      adc_rom[442] <= 4774;
      adc_rom[443] <= 4780;
      adc_rom[444] <= 4772;
      adc_rom[445] <= 4780;
      adc_rom[446] <= 4775;
      adc_rom[447] <= 4779;
      adc_rom[448] <= 4778;
      adc_rom[449] <= 4776;
      adc_rom[450] <= 4778;
      adc_rom[451] <= 4777;
      adc_rom[452] <= 4778;
      adc_rom[453] <= 4778;
      adc_rom[454] <= 4773;
      adc_rom[455] <= 4779;
      adc_rom[456] <= 4772;
      adc_rom[457] <= 4779;
      adc_rom[458] <= 4780;
      adc_rom[459] <= 4775;
      adc_rom[460] <= 4776;
      adc_rom[461] <= 4776;
      adc_rom[462] <= 4773;
      adc_rom[463] <= 4777;
      adc_rom[464] <= 4774;
      adc_rom[465] <= 4780;
      adc_rom[466] <= 4775;
      adc_rom[467] <= 4779;
      adc_rom[468] <= 4779;
      adc_rom[469] <= 4778;
      adc_rom[470] <= 4780;
      adc_rom[471] <= 4773;
      adc_rom[472] <= 4778;
      adc_rom[473] <= 4779;
      adc_rom[474] <= 4772;
      adc_rom[475] <= 4780;
      adc_rom[476] <= 4778;
      adc_rom[477] <= 4774;
      adc_rom[478] <= 4778;
      adc_rom[479] <= 4771;
      adc_rom[480] <= 4776;
      adc_rom[481] <= 4776;
      adc_rom[482] <= 4775;
      adc_rom[483] <= 4775;
      adc_rom[484] <= 4773;
      adc_rom[485] <= 4781;
      adc_rom[486] <= 4772;
      adc_rom[487] <= 4779;
      adc_rom[488] <= 4779;
      adc_rom[489] <= 4772;
      adc_rom[490] <= 4779;
      adc_rom[491] <= 4776;
      adc_rom[492] <= 4780;
      adc_rom[493] <= 4779;
      adc_rom[494] <= 4774;
      adc_rom[495] <= 4778;
      adc_rom[496] <= 4776;
      adc_rom[497] <= 4774;
      adc_rom[498] <= 4780;
      adc_rom[499] <= 4778;
      adc_rom[500] <= 4782;
      adc_rom[501] <= 4779;
      adc_rom[502] <= 4773;
      adc_rom[503] <= 4781;
      adc_rom[504] <= 4774;
      adc_rom[505] <= 4783;
      adc_rom[506] <= 4778;
      adc_rom[507] <= 4775;
      adc_rom[508] <= 4775;
      adc_rom[509] <= 4777;
      adc_rom[510] <= 4776;
      adc_rom[511] <= 4779;
      
   end
   
endmodule
